-- TestBench Template 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.std_logic_signed.all;
USE ieee.numeric_std.ALL;


  ENTITY testbench IS
  END testbench;

  ARCHITECTURE behavior OF testbench IS 



	--SIGNAL clk20us :  std_logic ;

   signal clk : std_logic := '0' ;
   signal input_I : signed(7 downto 0) := "00000000";
	signal input_Q : signed(7 downto 0) := "00000000";
   signal newValue : std_logic ;
 
	signal done_symbol : std_logic;

	signal output_value : std_logic;
	
	signal ascii_byte:  std_logic_vector(6 downto 0);
	

--constant clk20us_period : time := 20 us;         -- 0.2Mhz clk32 
constant clk_period : time := 10 ns;


BEGIN

	-- Instantiate the Unit Under Test (UUT)
	uut: entity work.top_counter PORT MAP(
		--clk20us => clk20us,
		clk  => clk ,
		input_I => input_I ,
	   input_Q => input_Q ,
	   newValue => newValue,
	   done => done_symbol,
		output_value => output_value,
		ascii_byte => ascii_byte);

   -- Clock process definitions
 --  clk20us_process :process
  -- begin
	--	clk20us <= '1';
	--	wait for clk20us_period/2;
	--	clk20us <= '0';
	--	wait for clk20us_period/2;
  -- end process;


 clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
	
	
	
	
	
	newValue_process :process
   begin
		newValue <= '0';
		wait for 19990 ns;
		newValue <= '1';
		wait for 10 ns;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;
		--WARNING: stops being accurate after 13 ms (MATLAB time) or 1.3 ms (VHDL time)
		
 
		input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
  input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00010000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 
		
		
		
 end process;




END;








