--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   22:16:58 05/07/2020
-- Design Name:   
-- Module Name:   D:/ise/ise_crack/code/testnco/testbetch.vhd
-- Project Name:  testnco
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: testnc
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_signed.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY testbetch IS
END testbetch;
 
ARCHITECTURE behavior OF testbetch IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT testnc
    PORT(
         rst : IN  std_logic;
         clk : IN  std_logic;
         clk_10ns : IN  std_logic;
			ena : in std_logic;
			
         input_signal : IN  std_logic_vector (7 downto 0);
       
			newValue : in std_logic ;
			
         sine_out : OUT  std_logic_vector(7 downto 0);
         cosine_out : OUT std_logic_vector (7 downto 0);
			
         df : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal rst : std_logic := '1';
   signal clk : std_logic := '0';
   signal clk_10ns : std_logic := '0';
	signal ena : std_logic := '1';
	
	
  -- signal input_I : signed (7 downto 0) := (others => '0');
  -- signal input_Q : signed (7 downto 0) := (others => '0');
  
   signal input_signal : std_logic_vector (7 downto 0) := (others => '0');
	
   signal newValue : std_logic := '0';

 	--Outputs
   signal sine_out : std_logic_vector(7 downto 0);
   signal cosine_out : std_logic_vector (7 downto 0);
	
   signal df : std_logic_vector(15 downto 0);

   -- Clock period definitions
   constant clk_period : time := 20 us;
	
   constant clk_10ns_period : time := 10 ns;
	
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: testnc PORT MAP (
          rst => rst,
          clk => clk,
			 ena => ena,
          clk_10ns => clk_10ns,
          --input_I => input_I,
         -- input_Q => input_Q,
			 input_signal => input_signal ,
          newValue => newValue,
          sine_out => sine_out ,
          cosine_out => cosine_out ,
          df => df
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   clk_10ns_process :process
   begin
		clk_10ns <= '0';
		wait for clk_10ns_period/2;
		clk_10ns <= '1';
		wait for clk_10ns_period/2;
   end process;
 


	newValue_process :process
   begin
		newValue <= '0';
		wait for 19990 ns;
		newValue <= '1';
		wait for 10 ns;
   end process;
 
 
 
 rst <= '0' after 100 ns;


 stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;
		--WARNING: stops being accurate after 13 ms (MATLAB time) or 1.3 ms (VHDL time)
	
input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00010000"; 
 wait for 20000 ns; 
 input_signal <= "11110000"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001111"; 
 wait for 20000 ns; 
 input_signal <= "11110001"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110010"; 
 wait for 20000 ns; 
 input_signal <= "00001110"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001101"; 
 wait for 20000 ns; 
 input_signal <= "11110011"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110100"; 
 wait for 20000 ns; 
 input_signal <= "00001100"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110101"; 
 wait for 20000 ns; 
 input_signal <= "00001011"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001010"; 
 wait for 20000 ns; 
 input_signal <= "11110110"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11110111"; 
 wait for 20000 ns; 
 input_signal <= "00001001"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00001000"; 
 wait for 20000 ns; 
 input_signal <= "11111000"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000000"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111111"; 
 wait for 20000 ns; 
 input_signal <= "00000001"; 
 wait for 20000 ns; 
 input_signal <= "11111110"; 
 wait for 20000 ns; 
 input_signal <= "00000010"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000011"; 
 wait for 20000 ns; 
 input_signal <= "11111101"; 
 wait for 20000 ns; 
 input_signal <= "00000100"; 
 wait for 20000 ns; 
 input_signal <= "11111100"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111011"; 
 wait for 20000 ns; 
 input_signal <= "00000101"; 
 wait for 20000 ns; 
 input_signal <= "11111010"; 
 wait for 20000 ns; 
 input_signal <= "00000110"; 
 wait for 20000 ns; 
 input_signal <= "11111001"; 
 wait for 20000 ns; 
 input_signal <= "00000111"; 
     
 end process;
END;

